----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01.05.2017 20:52:12
-- Design Name: 
-- Module Name: top - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity StaticPlaceholder is
    Port ( 
    
    NET_Left_X1Y5_out    : out std_logic_vector(215 downto 0);
    NET_Left_X1Y5_in     : in std_logic_vector(215 downto 0);
    NET_Right_X1Y5_out   : out std_logic_vector(215 downto 0);
    NET_Right_X1Y5_in    : in std_logic_vector(215 downto 0));
    
    
end StaticPlaceholder;

architecture Behavioral of StaticPlaceholder is

constant size : integer := 54;

attribute MARK_DEBUG : string;

-- START_DECLARATION
-- END_DECLARATION

signal NET_X1Y5_west        : std_logic_vector((size*4)-1 downto 0);
signal NET_X1Y5_east        : std_logic_vector((size*4)-1 downto 0);
--signal NET_Left_X1Y5_out    : std_logic_vector((size*4)-1 downto 0);
--signal NET_Left_X1Y5_in     : std_logic_vector((size*4)-1 downto 0);
--signal NET_Right_X1Y5_out   : std_logic_vector((size*4)-1 downto 0);
--signal NET_Right_X1Y5_in    : std_logic_vector((size*4)-1 downto 0);

attribute MARK_DEBUG of  NET_X1Y5_west :  signal is "TRUE";
attribute MARK_DEBUG of  NET_X1Y5_east :  signal is "TRUE";
attribute MARK_DEBUG of  NET_Left_X1Y5_out :  signal is "TRUE";
attribute MARK_DEBUG of  NET_Right_X1Y5_out :  signal is "TRUE";

begin
--# >>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>> 
--# [NET_Left_X1Y5_in(0)] G1 -> GQ  -> [NET_X1Y5_east(0)] EE4_E_BEG4 -> EE2_E_END4 -> IMUX_E36  G4 -> GQ  [NET_Right_X1Y5_out(0)]     EE2_E_END4 -> INT_NODE_IMUX_14_INT_OUT0 -> was_IMUX_E36_G4_
--# [NET_Left_X1Y5_in(1)] G2 -> GQ2 -> [NET_X1Y5_east(1)] EE4_E_BEG2 -> EE2_E_END2 -> IMUX_E3   F1 -> FQ2 [NET_Right_X1Y5_out(1)]    EE2_E_END2 -> INT_NODE_IMUX_4_INT_OUT1  -> was_IMUX_E3_F1_
--# [NET_Left_X1Y5_in(2)] H1 -> HQ  -> [NET_X1Y5_east(2)] EE4_E_BEG6 -> EE2_E_END6 -> IMUX_E14  G2 -> GQ2 [NET_Right_X1Y5_out(2)]    EE2_E_END6 -> INT_NODE_IMUX_23_INT_OUT0 -> was_IMUX_E14_G2_
--# [NET_Left_X1Y5_in(3)] F1 -> FQ2 -> [NET_X1Y5_east(3)] EE4_E_BEG0 -> EE2_E_END0 -> IMUX_E1   H1 -> HQ  [NET_Right_X1Y5_out(3)]    EE2_E_END0 -> INT_NODE_IMUX_11_INT_OUT0 -> was_IMUX_E1_H1_
--# the right LUT inputs leave us little choice G4, F1, G2, H1;  These are not allowed on the other side (left) (for the WW direction)

--# <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<
--# [NET_Left_X1Y5_out(0)] EQ 	<- IMUX_E40  E3 <- WW2_E_END7 <- WW4_E_BEG7 [NET_X1Y5_west(0)] <- EQ  <- E1  [NET_Right_X1Y5_in(0)]    WW2_E_END7 -> INT_NODE_IMUX_27_INT_OUT1 -> was_IMUX_E40_E3_   
--# [NET_Left_X1Y5_out(1)] EQ2	<- IMUX_E4   E2 <- WW2_E_END1 <- WW4_E_BEG1 [NET_X1Y5_west(1)] <- EQ2 <- E2  [NET_Right_X1Y5_in(1)]    WW2_E_END1 -> INT_NODE_IMUX_1_INT_OUT0 -> was_IMUX_E4_E2_
--# [NET_Left_X1Y5_out(2)] HQ2	<- IMUX_E33  H3 <- WW2_E_END3 <- WW4_E_BEG3 [NET_X1Y5_west(2)] <- HQ2 <- H2  [NET_Right_X1Y5_in(2)]    WW2_E_END3 -> INT_NODE_IMUX_10_INT_OUT0 -> was_IMUX_E33_H3_
--# [NET_Left_X1Y5_out(3)] FQ 	<- IMUX_E41  F3 <- WW2_E_END5 <- WW4_E_BEG5 [NET_X1Y5_west(3)] <- FQ  <- F2  [NET_Right_X1Y5_in(3)]    WW2_E_END5 -> INT_NODE_IMUX_19_INT_OUT0 -> was_IMUX_E41_F3_    WW2_E_END5 -> INT_NODE_IMUX_18_INT_OUT0 -> was_IMUX_E43_F5_
--# the left LUT inputs leave us little choice E3, E2, H3, F3;  These are not allowed on the other side (right) (for the EE direction)

-- START_BODY

INST_Left_X1Y5_E6LUT_0 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(0), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(1), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(1), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(0), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_0 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(3), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(3), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(3), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(3), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_0 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(0), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(1), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(0), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(1), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_0 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(2), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(2), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(2), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(2), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_0 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(0), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(1), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(0), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(1), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_0 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(3), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(1), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(1), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(3), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_0 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(0), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(2), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(2), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(0), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_0 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(3), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(2), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(3), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(2), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_1 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(4), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(5), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(5), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(4), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_1 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(7), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(7), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(7), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(7), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_1 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(4), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(5), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(4), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(5), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_1 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(6), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(6), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(6), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(6), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_1 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(4), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(5), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(4), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(5), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_1 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(7), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(5), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(5), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(7), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_1 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(4), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(6), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(6), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(4), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_1 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(7), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(6), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(7), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(6), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_2 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(8), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(9), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(9), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(8), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_2 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(11), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(11), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(11), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(11), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_2 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(8), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(9), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(8), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(9), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_2 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(10), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(10), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(10), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(10), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_2 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(8), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(9), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(8), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(9), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_2 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(11), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(9), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(9), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(11), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_2 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(8), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(10), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(10), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(8), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_2 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(11), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(10), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(11), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(10), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_3 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(12), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(13), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(13), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(12), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_3 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(15), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(15), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(15), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(15), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_3 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(12), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(13), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(12), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(13), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_3 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(14), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(14), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(14), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(14), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_3 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(12), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(13), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(12), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(13), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_3 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(15), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(13), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(13), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(15), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_3 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(12), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(14), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(14), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(12), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_3 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(15), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(14), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(15), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(14), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_4 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(16), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(17), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(17), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(16), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_4 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(19), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(19), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(19), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(19), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_4 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(16), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(17), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(16), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(17), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_4 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(18), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(18), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(18), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(18), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_4 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(16), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(17), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(16), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(17), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_4 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(19), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(17), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(17), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(19), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_4 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(16), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(18), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(18), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(16), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_4 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(19), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(18), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(19), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(18), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_5 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(20), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(21), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(21), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(20), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_5 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(23), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(23), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(23), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(23), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_5 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(20), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(21), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(20), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(21), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_5 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(22), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(22), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(22), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(22), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_5 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(20), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(21), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(20), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(21), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_5 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(23), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(21), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(21), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(23), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_5 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(20), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(22), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(22), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(20), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_5 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(23), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(22), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(23), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(22), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_6 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(24), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(25), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(25), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(24), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_6 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(27), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(27), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(27), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(27), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_6 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(24), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(25), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(24), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(25), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_6 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(26), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(26), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(26), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(26), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_6 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(24), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(25), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(24), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(25), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_6 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(27), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(25), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(25), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(27), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_6 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(24), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(26), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(26), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(24), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_6 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(27), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(26), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(27), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(26), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_7 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(28), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(29), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(29), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(28), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_7 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(31), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(31), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(31), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(31), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_7 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(28), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(29), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(28), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(29), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_7 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(30), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(30), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(30), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(30), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_7 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(28), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(29), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(28), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(29), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_7 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(31), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(29), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(29), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(31), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_7 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(28), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(30), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(30), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(28), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_7 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(31), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(30), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(31), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(30), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_8 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(32), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(33), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(33), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(32), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_8 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(35), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(35), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(35), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(35), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_8 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(32), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(33), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(32), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(33), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_8 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(34), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(34), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(34), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(34), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_8 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(32), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(33), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(32), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(33), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_8 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(35), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(33), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(33), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(35), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_8 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(32), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(34), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(34), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(32), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_8 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(35), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(34), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(35), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(34), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_9 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(36), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(37), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(37), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(36), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_9 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(39), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(39), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(39), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(39), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_9 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(36), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(37), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(36), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(37), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_9 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(38), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(38), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(38), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(38), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_9 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(36), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(37), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(36), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(37), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_9 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(39), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(37), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(37), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(39), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_9 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(36), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(38), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(38), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(36), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_9 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(39), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(38), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(39), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(38), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_10 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(40), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(41), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(41), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(40), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_10 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(43), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(43), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(43), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(43), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_10 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(40), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(41), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(40), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(41), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_10 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(42), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(42), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(42), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(42), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_10 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(40), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(41), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(40), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(41), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_10 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(43), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(41), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(41), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(43), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_10 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(40), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(42), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(42), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(40), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_10 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(43), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(42), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(43), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(42), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_11 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(44), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(45), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(45), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(44), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_11 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(47), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(47), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(47), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(47), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_11 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(44), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(45), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(44), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(45), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_11 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(46), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(46), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(46), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(46), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_11 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(44), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(45), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(44), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(45), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_11 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(47), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(45), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(45), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(47), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_11 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(44), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(46), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(46), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(44), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_11 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(47), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(46), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(47), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(46), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_12 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(48), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(49), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(49), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(48), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_12 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(51), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(51), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(51), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(51), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_12 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(48), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(49), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(48), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(49), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_12 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(50), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(50), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(50), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(50), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_12 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(48), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(49), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(48), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(49), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_12 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(51), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(49), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(49), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(51), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_12 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(48), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(50), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(50), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(48), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_12 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(51), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(50), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(51), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(50), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_13 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(52), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(53), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(53), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(52), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_13 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(55), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(55), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(55), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(55), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_13 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(52), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(53), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(52), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(53), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_13 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(54), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(54), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(54), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(54), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_13 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(52), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(53), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(52), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(53), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_13 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(55), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(53), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(53), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(55), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_13 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(52), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(54), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(54), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(52), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_13 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(55), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(54), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(55), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(54), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_14 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(56), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(57), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(57), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(56), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_14 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(59), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(59), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(59), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(59), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_14 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(56), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(57), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(56), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(57), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_14 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(58), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(58), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(58), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(58), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_14 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(56), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(57), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(56), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(57), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_14 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(59), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(57), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(57), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(59), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_14 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(56), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(58), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(58), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(56), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_14 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(59), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(58), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(59), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(58), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_15 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(60), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(61), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(61), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(60), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_15 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(63), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(63), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(63), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(63), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_15 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(60), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(61), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(60), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(61), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_15 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(62), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(62), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(62), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(62), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_15 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(60), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(61), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(60), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(61), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_15 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(63), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(61), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(61), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(63), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_15 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(60), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(62), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(62), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(60), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_15 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(63), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(62), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(63), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(62), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_16 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(64), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(65), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(65), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(64), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_16 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(67), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(67), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(67), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(67), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_16 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(64), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(65), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(64), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(65), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_16 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(66), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(66), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(66), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(66), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_16 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(64), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(65), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(64), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(65), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_16 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(67), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(65), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(65), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(67), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_16 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(64), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(66), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(66), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(64), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_16 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(67), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(66), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(67), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(66), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_17 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(68), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(69), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(69), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(68), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_17 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(71), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(71), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(71), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(71), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_17 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(68), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(69), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(68), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(69), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_17 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(70), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(70), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(70), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(70), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_17 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(68), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(69), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(68), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(69), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_17 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(71), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(69), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(69), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(71), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_17 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(68), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(70), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(70), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(68), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_17 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(71), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(70), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(71), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(70), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_18 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(72), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(73), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(73), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(72), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_18 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(75), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(75), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(75), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(75), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_18 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(72), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(73), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(72), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(73), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_18 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(74), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(74), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(74), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(74), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_18 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(72), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(73), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(72), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(73), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_18 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(75), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(73), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(73), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(75), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_18 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(72), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(74), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(74), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(72), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_18 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(75), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(74), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(75), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(74), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_19 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(76), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(77), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(77), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(76), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_19 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(79), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(79), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(79), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(79), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_19 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(76), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(77), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(76), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(77), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_19 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(78), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(78), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(78), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(78), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_19 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(76), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(77), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(76), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(77), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_19 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(79), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(77), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(77), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(79), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_19 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(76), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(78), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(78), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(76), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_19 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(79), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(78), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(79), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(78), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_20 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(80), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(81), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(81), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(80), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_20 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(83), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(83), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(83), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(83), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_20 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(80), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(81), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(80), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(81), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_20 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(82), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(82), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(82), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(82), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_20 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(80), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(81), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(80), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(81), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_20 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(83), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(81), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(81), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(83), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_20 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(80), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(82), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(82), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(80), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_20 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(83), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(82), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(83), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(82), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_21 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(84), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(85), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(85), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(84), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_21 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(87), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(87), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(87), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(87), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_21 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(84), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(85), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(84), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(85), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_21 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(86), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(86), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(86), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(86), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_21 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(84), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(85), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(84), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(85), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_21 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(87), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(85), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(85), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(87), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_21 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(84), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(86), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(86), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(84), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_21 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(87), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(86), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(87), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(86), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_22 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(88), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(89), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(89), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(88), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_22 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(91), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(91), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(91), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(91), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_22 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(88), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(89), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(88), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(89), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_22 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(90), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(90), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(90), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(90), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_22 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(88), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(89), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(88), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(89), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_22 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(91), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(89), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(89), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(91), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_22 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(88), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(90), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(90), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(88), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_22 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(91), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(90), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(91), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(90), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_23 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(92), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(93), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(93), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(92), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_23 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(95), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(95), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(95), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(95), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_23 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(92), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(93), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(92), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(93), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_23 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(94), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(94), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(94), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(94), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_23 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(92), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(93), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(92), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(93), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_23 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(95), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(93), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(93), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(95), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_23 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(92), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(94), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(94), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(92), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_23 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(95), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(94), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(95), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(94), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_24 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(96), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(97), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(97), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(96), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_24 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(99), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(99), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(99), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(99), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_24 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(96), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(97), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(96), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(97), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_24 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(98), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(98), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(98), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(98), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_24 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(96), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(97), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(96), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(97), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_24 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(99), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(97), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(97), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(99), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_24 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(96), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(98), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(98), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(96), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_24 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(99), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(98), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(99), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(98), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_25 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(100), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(101), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(101), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(100), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_25 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(103), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(103), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(103), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(103), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_25 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(100), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(101), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(100), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(101), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_25 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(102), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(102), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(102), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(102), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_25 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(100), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(101), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(100), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(101), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_25 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(103), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(101), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(101), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(103), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_25 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(100), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(102), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(102), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(100), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_25 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(103), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(102), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(103), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(102), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_26 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(104), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(105), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(105), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(104), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_26 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(107), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(107), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(107), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(107), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_26 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(104), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(105), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(104), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(105), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_26 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(106), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(106), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(106), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(106), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_26 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(104), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(105), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(104), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(105), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_26 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(107), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(105), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(105), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(107), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_26 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(104), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(106), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(106), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(104), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_26 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(107), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(106), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(107), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(106), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_27 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(108), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(109), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(109), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(108), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_27 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(111), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(111), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(111), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(111), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_27 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(108), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(109), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(108), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(109), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_27 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(110), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(110), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(110), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(110), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_27 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(108), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(109), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(108), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(109), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_27 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(111), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(109), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(109), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(111), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_27 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(108), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(110), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(110), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(108), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_27 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(111), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(110), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(111), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(110), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_28 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(112), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(113), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(113), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(112), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_28 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(115), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(115), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(115), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(115), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_28 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(112), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(113), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(112), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(113), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_28 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(114), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(114), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(114), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(114), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_28 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(112), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(113), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(112), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(113), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_28 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(115), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(113), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(113), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(115), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_28 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(112), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(114), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(114), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(112), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_28 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(115), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(114), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(115), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(114), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_29 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(116), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(117), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(117), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(116), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_29 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(119), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(119), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(119), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(119), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_29 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(116), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(117), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(116), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(117), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_29 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(118), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(118), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(118), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(118), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_29 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(116), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(117), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(116), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(117), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_29 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(119), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(117), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(117), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(119), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_29 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(116), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(118), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(118), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(116), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_29 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(119), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(118), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(119), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(118), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_30 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(120), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(121), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(121), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(120), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_30 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(123), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(123), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(123), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(123), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_30 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(120), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(121), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(120), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(121), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_30 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(122), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(122), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(122), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(122), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_30 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(120), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(121), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(120), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(121), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_30 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(123), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(121), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(121), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(123), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_30 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(120), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(122), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(122), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(120), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_30 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(123), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(122), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(123), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(122), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_31 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(124), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(125), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(125), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(124), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_31 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(127), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(127), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(127), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(127), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_31 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(124), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(125), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(124), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(125), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_31 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(126), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(126), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(126), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(126), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_31 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(124), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(125), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(124), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(125), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_31 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(127), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(125), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(125), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(127), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_31 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(124), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(126), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(126), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(124), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_31 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(127), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(126), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(127), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(126), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_32 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(128), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(129), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(129), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(128), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_32 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(131), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(131), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(131), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(131), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_32 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(128), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(129), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(128), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(129), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_32 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(130), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(130), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(130), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(130), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_32 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(128), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(129), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(128), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(129), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_32 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(131), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(129), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(129), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(131), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_32 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(128), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(130), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(130), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(128), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_32 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(131), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(130), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(131), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(130), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_33 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(132), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(133), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(133), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(132), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_33 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(135), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(135), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(135), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(135), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_33 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(132), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(133), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(132), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(133), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_33 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(134), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(134), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(134), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(134), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_33 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(132), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(133), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(132), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(133), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_33 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(135), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(133), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(133), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(135), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_33 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(132), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(134), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(134), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(132), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_33 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(135), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(134), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(135), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(134), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_34 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(136), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(137), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(137), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(136), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_34 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(139), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(139), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(139), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(139), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_34 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(136), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(137), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(136), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(137), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_34 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(138), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(138), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(138), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(138), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_34 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(136), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(137), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(136), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(137), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_34 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(139), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(137), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(137), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(139), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_34 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(136), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(138), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(138), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(136), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_34 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(139), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(138), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(139), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(138), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_35 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(140), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(141), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(141), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(140), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_35 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(143), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(143), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(143), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(143), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_35 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(140), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(141), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(140), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(141), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_35 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(142), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(142), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(142), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(142), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_35 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(140), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(141), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(140), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(141), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_35 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(143), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(141), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(141), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(143), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_35 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(140), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(142), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(142), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(140), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_35 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(143), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(142), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(143), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(142), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_36 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(144), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(145), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(145), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(144), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_36 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(147), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(147), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(147), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(147), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_36 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(144), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(145), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(144), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(145), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_36 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(146), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(146), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(146), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(146), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_36 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(144), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(145), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(144), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(145), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_36 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(147), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(145), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(145), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(147), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_36 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(144), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(146), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(146), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(144), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_36 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(147), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(146), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(147), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(146), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_37 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(148), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(149), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(149), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(148), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_37 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(151), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(151), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(151), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(151), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_37 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(148), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(149), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(148), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(149), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_37 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(150), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(150), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(150), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(150), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_37 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(148), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(149), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(148), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(149), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_37 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(151), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(149), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(149), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(151), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_37 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(148), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(150), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(150), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(148), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_37 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(151), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(150), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(151), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(150), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_38 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(152), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(153), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(153), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(152), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_38 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(155), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(155), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(155), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(155), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_38 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(152), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(153), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(152), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(153), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_38 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(154), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(154), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(154), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(154), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_38 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(152), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(153), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(152), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(153), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_38 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(155), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(153), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(153), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(155), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_38 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(152), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(154), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(154), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(152), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_38 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(155), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(154), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(155), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(154), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_39 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(156), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(157), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(157), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(156), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_39 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(159), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(159), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(159), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(159), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_39 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(156), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(157), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(156), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(157), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_39 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(158), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(158), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(158), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(158), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_39 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(156), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(157), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(156), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(157), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_39 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(159), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(157), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(157), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(159), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_39 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(156), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(158), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(158), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(156), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_39 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(159), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(158), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(159), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(158), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_40 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(160), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(161), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(161), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(160), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_40 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(163), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(163), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(163), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(163), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_40 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(160), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(161), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(160), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(161), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_40 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(162), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(162), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(162), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(162), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_40 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(160), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(161), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(160), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(161), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_40 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(163), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(161), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(161), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(163), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_40 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(160), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(162), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(162), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(160), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_40 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(163), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(162), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(163), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(162), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_41 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(164), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(165), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(165), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(164), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_41 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(167), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(167), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(167), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(167), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_41 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(164), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(165), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(164), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(165), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_41 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(166), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(166), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(166), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(166), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_41 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(164), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(165), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(164), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(165), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_41 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(167), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(165), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(165), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(167), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_41 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(164), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(166), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(166), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(164), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_41 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(167), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(166), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(167), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(166), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_42 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(168), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(169), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(169), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(168), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_42 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(171), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(171), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(171), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(171), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_42 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(168), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(169), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(168), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(169), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_42 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(170), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(170), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(170), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(170), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_42 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(168), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(169), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(168), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(169), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_42 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(171), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(169), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(169), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(171), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_42 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(168), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(170), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(170), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(168), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_42 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(171), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(170), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(171), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(170), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_43 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(172), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(173), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(173), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(172), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_43 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(175), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(175), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(175), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(175), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_43 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(172), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(173), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(172), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(173), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_43 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(174), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(174), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(174), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(174), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_43 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(172), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(173), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(172), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(173), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_43 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(175), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(173), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(173), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(175), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_43 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(172), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(174), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(174), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(172), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_43 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(175), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(174), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(175), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(174), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_44 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(176), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(177), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(177), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(176), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_44 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(179), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(179), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(179), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(179), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_44 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(176), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(177), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(176), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(177), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_44 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(178), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(178), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(178), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(178), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_44 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(176), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(177), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(176), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(177), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_44 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(179), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(177), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(177), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(179), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_44 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(176), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(178), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(178), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(176), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_44 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(179), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(178), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(179), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(178), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_45 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(180), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(181), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(181), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(180), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_45 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(183), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(183), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(183), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(183), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_45 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(180), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(181), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(180), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(181), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_45 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(182), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(182), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(182), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(182), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_45 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(180), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(181), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(180), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(181), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_45 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(183), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(181), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(181), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(183), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_45 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(180), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(182), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(182), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(180), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_45 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(183), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(182), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(183), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(182), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_46 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(184), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(185), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(185), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(184), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_46 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(187), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(187), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(187), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(187), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_46 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(184), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(185), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(184), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(185), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_46 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(186), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(186), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(186), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(186), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_46 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(184), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(185), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(184), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(185), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_46 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(187), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(185), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(185), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(187), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_46 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(184), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(186), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(186), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(184), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_46 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(187), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(186), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(187), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(186), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_47 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(188), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(189), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(189), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(188), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_47 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(191), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(191), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(191), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(191), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_47 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(188), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(189), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(188), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(189), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_47 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(190), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(190), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(190), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(190), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_47 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(188), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(189), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(188), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(189), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_47 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(191), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(189), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(189), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(191), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_47 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(188), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(190), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(190), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(188), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_47 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(191), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(190), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(191), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(190), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_48 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(192), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(193), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(193), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(192), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_48 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(195), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(195), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(195), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(195), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_48 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(192), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(193), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(192), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(193), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_48 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(194), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(194), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(194), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(194), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_48 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(192), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(193), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(192), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(193), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_48 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(195), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(193), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(193), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(195), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_48 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(192), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(194), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(194), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(192), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_48 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(195), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(194), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(195), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(194), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_49 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(196), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(197), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(197), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(196), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_49 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(199), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(199), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(199), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(199), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_49 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(196), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(197), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(196), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(197), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_49 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(198), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(198), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(198), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(198), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_49 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(196), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(197), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(196), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(197), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_49 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(199), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(197), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(197), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(199), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_49 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(196), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(198), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(198), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(196), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_49 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(199), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(198), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(199), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(198), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_50 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(200), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(201), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(201), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(200), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_50 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(203), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(203), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(203), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(203), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_50 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(200), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(201), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(200), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(201), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_50 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(202), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(202), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(202), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(202), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_50 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(200), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(201), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(200), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(201), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_50 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(203), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(201), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(201), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(203), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_50 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(200), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(202), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(202), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(200), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_50 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(203), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(202), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(203), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(202), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_51 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(204), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(205), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(205), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(204), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_51 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(207), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(207), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(207), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(207), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_51 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(204), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(205), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(204), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(205), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_51 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(206), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(206), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(206), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(206), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_51 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(204), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(205), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(204), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(205), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_51 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(207), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(205), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(205), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(207), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_51 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(204), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(206), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(206), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(204), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_51 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(207), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(206), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(207), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(206), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_52 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(208), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(209), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(209), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(208), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_52 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(211), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(211), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(211), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(211), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_52 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(208), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(209), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(208), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(209), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_52 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(210), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(210), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(210), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(210), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_52 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(208), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(209), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(208), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(209), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_52 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(211), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(209), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(209), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(211), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_52 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(208), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(210), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(210), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(208), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_52 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(211), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(210), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(211), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(210), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );




INST_Left_X1Y5_E6LUT_53 : LUT6_2
generic map (
INIT => X"F0F0F0F0CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(212), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(213), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- E1 LUT input (1-bit) 
		   I1 => NET_X1Y5_west(213), -- E2 LUT input (1-bit)
           I2 => NET_X1Y5_west(212), -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Left_X1Y5_D6LUT_53 : LUT6_2
generic map (
INIT => X"F0F0F0F0AAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_Left_X1Y5_out(215), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(215), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(215), -- F1 LUT input (1-bit) 
		   I1 => '1', -- F2 LUT input (1-bit)
           I2 => NET_X1Y5_west(215), -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Left_X1Y5_G6LUT_53 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(212), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_east(213), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(212), -- G1 LUT input (1-bit) 
		   I1 => NET_Left_X1Y5_in(213), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => '1', -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Left_X1Y5_C6LUT_53 : LUT6_2
generic map (
INIT => X"AAAAAAAAF0F0F0F0") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_east(214), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Left_X1Y5_out(214), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Left_X1Y5_in(214), -- H1 LUT input (1-bit) 
		   I1 => '1', -- H2 LUT input (1-bit)
           I2 => NET_X1Y5_west(214), -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );
 
          
 
          
-- Right side
INST_Right_X1Y5_E6LUT_53 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(212), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(213), -- to Q2 5-LUT output (1-bit)
           I0 => NET_Right_X1Y5_in(212), -- E1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(213), -- E2 LUT input (1-bit)
           I2 => '1', -- E3 LUT input (1-bit)
           I3 => '1', -- E4 LUT input (1-bit)
           I4 => '1', -- E5 LUT input (1-bit)
           I5 => '1'  -- E6 LUT input (1-bit)
         );

INST_Right_X1Y5_D6LUT_53 : LUT6_2
generic map (
INIT => X"CCCCCCCCAAAAAAAA") -- Specify LUT Contents 
port map ( O6 => NET_X1Y5_west(215), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(213), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(213), -- F1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(215), -- F2 LUT input (1-bit)
           I2 => '1', -- F3 LUT input (1-bit)
           I3 => '1', -- F4 LUT input (1-bit)
           I4 => '1', -- F5 LUT input (1-bit)
           I5 => '1'  -- D6 LUT input (1-bit)
         );

INST_Right_X1Y5_G6LUT_53 : LUT6_2
generic map (
INIT => X"FF00FF00CCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(212), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_Right_X1Y5_out(214), -- to Q2 5-LUT output (1-bit)
           I0 => '1', -- G1 LUT input (1-bit) 
		   I1 => NET_X1Y5_east(214), -- G2 LUT input (1-bit)
           I2 => '1', -- G3 LUT input (1-bit)
           I3 => NET_X1Y5_east(212), -- G4 LUT input (1-bit)
           I4 => '1', -- G5 LUT input (1-bit)
           I5 => '1'  -- G6 LUT input (1-bit)
         );

INST_Right_X1Y5_C6LUT_53 : LUT6_2
generic map (
INIT => X"AAAAAAAACCCCCCCC") -- Specify LUT Contents 
port map ( O6 => NET_Right_X1Y5_out(215), -- to Q 6/5-LUT output (1-bit)
           O5 => NET_X1Y5_west(214), -- to Q2 5-LUT output (1-bit)
           I0 => NET_X1Y5_east(215), -- H1 LUT input (1-bit) 
		   I1 => NET_Right_X1Y5_in(214), -- H2 LUT input (1-bit)
           I2 => '1', -- H3 LUT input (1-bit)
           I3 => '1', -- H4 LUT input (1-bit)
           I4 => '1', -- H5 LUT input (1-bit)
           I5 => '1'  -- C6 LUT input (1-bit)
         );



-- END_BODY

end Behavioral;
